// Parameters for DUT and OVL checker

// number of data bits
// WIDTH = B

`define B 8
`define WIDTH 8

// depth or number of adress bits
// DEPTH = 2**W

`define W 5
`define DEPTH 32

// clock period

`define PERIOD 100
